`timescale 1ns/1ns
module MUX_8_1_tb;
	reg [15:0]A0;
	reg [15:0]A1;
	reg [15:0]A2;
	reg [15:0]A3;
	reg [15:0]A4;
	reg [15:0]A5;
	reg [15:0]A6;
	reg [15:0]A7;
	reg [2:0]S;
	wire [15:0]O;

	MUX_8_1 muxTest(.a0(A0),.a1(A1),.a2(A2),.a3(A3),.a4(A4),.a5(A5),.a6(A6),.a7(A7),.s(S),.o(O));

	initial begin
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b000;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b001;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b010;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b011;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b100;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b101;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b110;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;S=3'b111;
	end
	initial begin
		$dumpfile("MUX_8_1.vcd");
		$dumpvars;
	end
endmodule
