`timescale 1ns/1ns
module MUX_16_1_tb;
	reg [15:0]A0;
	reg [15:0]A1;
	reg [15:0]A2;
	reg [15:0]A3;
	reg [15:0]A4;
	reg [15:0]A5;
	reg [15:0]A6;
	reg [15:0]A7;
	reg [15:0]A8;
	reg [15:0]A9;
	reg [15:0]A10;
	reg [15:0]A11;
	reg [15:0]A12;
	reg [15:0]A13;
	reg [15:0]A14;
	reg [15:0]A15;
	reg [3:0]S;
	wire [15:0]O;

	MUX_16_1 muxTest(.a0(A0),.a1(A1),.a2(A2),.a3(A3),.a4(A4),.a5(A5),.a6(A6),.a7(A7),.a8(A8),.a9(A9),.a10(A10),.a11(A11),.a12(A12),.a13(A13),.a14(A14),.a15(A15),.s(S),.o(O));

	initial begin
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0000;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0001;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0010;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0011;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0100;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0101;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0110;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b0111;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1000;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1001;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1010;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1011;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1100;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1101;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1110;
		#1
		A0=4'b0001;A1=4'b0010;A2=4'b0011;A3=4'b0100;A4=4'b0101;A5=4'b0110;A6=4'b0111;A7=4'b1000;A8=4'b1001;A9=4'b1010;A10=4'b1011;A11=4'b1100;A12=4'b1101;A13=4'b1110;A14=4'b1111;A15=4'b0000;S=4'b1111;
	end
	initial begin
		$dumpfile("MUX_16_1.vcd");
		$dumpvars;
	end
endmodule
